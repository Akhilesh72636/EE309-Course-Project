library ieee;
use ieee.std_logic_1164.all;

entity registers_file is 
    port(
        
        A1 : in std_logic_vector(2 downto 0); -- to store register adress 
        A2 : in std_logic_vector(2 downto 0); -- to store register adress 
        A3 : in std_logic_vector(2 downto 0); -- to store register adress
		  
        -- input data
        Din : in std_logic_vector(15 downto 0);-- input data to store in register
		  R0in : in std_logic_vector(15 downto 0);
		  WR_ER0: in std_logic;
        WR_E : in std_logic; -- write enable
        reset : in std_logic; -- reset input
        clk : in std_logic; --clock
        --output data
        D1 : out std_logic_vector(15 downto 0); -- data output 1
        D2 : out std_logic_vector(15 downto 0); -- data output 2
        R0_PC : out std_logic_vector(15 downto 0)  -- value of R7 as pc

    );
end entity;

architecture inside of registers_file is    
    signal R0 : std_logic_vector(15 downto 0) ;
    signal R1 : std_logic_vector(15 downto 0) ;
    signal R2 : std_logic_vector(15 downto 0) ;
    signal R3 : std_logic_vector(15 downto 0);
    signal R4 : std_logic_vector(15 downto 0) ;
    signal R5 : std_logic_vector(15 downto 0);
    signal R6 : std_logic_vector(15 downto 0);
    signal R7 : std_logic_vector(15 downto 0);
	 
	
	begin
    
    write_process: process(A3,WR_E,clk,reset,WR_ER0,R0in) --writing to register when write_enable is set
    begin
	 
	    if(reset = '1') then             --initiating all values of Rrgister to "0"
            R0 <= "0000000000000000";
            R1 <= "0000000000000000";
            R2 <= "0000000000000000";
            R3 <= "0000000000000000";
            R4 <= "0000000000000000";
            R5 <= "0000000000000000";
            R6 <= "0000000000000000";
            R7 <= "0000000000000000";
				
elsif (clk'event and clk = '1') then  --writing data in registers 
   if(WR_ER0 = '1') then
     --writing  in register  R0
                    R0 <= R0in;
end if;						  
	if(WR_E = '1') then
				
                if(A3 = "000") then     --writing  in register  R0
                    R0 <= Din;
                
                elsif(A3 = "001") then
                    R1 <= Din;
						  
                elsif(A3 = "010") then
                    R2 <= Din;
						  
                elsif(A3 = "011") then
                    R3 <= Din;

                elsif(A3 = "100") then
                    R4 <= Din;

                elsif(A3 = "101") then
                    R5 <= Din;
	
                elsif(A3 = "110") then
                    R6 <= Din;
 		 
                elsif(A3 = "111") then
                    R7 <= Din;
                end if;
    end if;
end if;
end process write_process;
	 
	
read_process: process(A1,A2) -- to read data from registers

begin
        
		
		
            if(A1 = "000")    then  -- to read data from registers to Data output D1
                D1 <= R0;

            elsif(A1 = "001") then
                D1 <= R1;
 
            elsif(A1 = "010") then
                D1 <= R2;
     
            elsif(A1 = "011") then
                D1 <= R3;
         
            elsif(A1 = "100") then
                D1 <= R4;
          
            elsif(A1 = "101") then
                D1 <= R5;
    
            elsif(A1 = "110") then
                D1 <= R6;
       
            elsif(A1 = "111") then
                D1 <= R7;
            end if;
				
           
            if(A2 = "000")    then     -- to read data from registers to Data output D1
                D2 <= R0;
            
            elsif(A2 = "001") then
                D2 <= R1;
            
            elsif(A2 = "010") then
                D2 <= R2;
          
            elsif(A2 = "011") then
                D2 <= R3;
          
            elsif(A2 = "100") then
                D2 <= R4;
          
            elsif(A2 = "101") then
                D2 <= R5;
            
            elsif(A2 = "110") then
                D2 <= R6;
        
            elsif(A2 = "111") then
                D2 <= R7;
            end if;    
  
      
    end process read_process;

    R0_PC <= R0;
end inside;