library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity EXMM_Reg is
	port (
	     clk: in std_logic;
        PCin : IN STD_LOGIC_VECTOR(15 downto 0);     ---------input 
		  WR_E: in std_logic;                          -- enable input
        reset: in std_logic;
		  Iin : IN STD_LOGIC_VECTOR(15 downto 0);
         opcodein: in STD_LOGIC_VECTOR(3 downto 0); 
			
			aluCin : in STD_LOGIC_VECTOR(15 downto 0);
			
		   Immin : in STD_LOGIC_VECTOR(15 downto 0);
			aRAin : in STD_LOGIC_VECTOR(2 downto 0);
			---------------------------------------------------
		  PCout : out STD_LOGIC_VECTOR(15 downto 0); 
		  Iout : out STD_LOGIC_VECTOR(15 downto 0) ; ------------ output
		   opcode: OUT STD_LOGIC_VECTOR(3 downto 0); 
			aluCout : out STD_LOGIC_VECTOR(15 downto 0);
			tellin:in std_logic;
			tellout:in std_logic;
			aRAout : out STD_LOGIC_VECTOR(2 downto 0);
		
		   Imm : OUT STD_LOGIC_VECTOR(15 downto 0));
end EXMM_Reg;


architecture behave of EXMM_Reg is
  begin 
  
    process(Iin,clk,PCin,reset,WR_E,opcodein,aluCin ,Immin,aRAin ,tellin ) is
	  variable T1, compvalue,One: STD_LOGIC_VECTOR(15 downto 0);
      begin
		if (clk'event and clk = '1') then
		  
		 if(reset='1') then
               Iout  <="----------------";
               PCout <="----------------"  ;
					opcode<="----";
			      aluCout<="----------------"; 
		         Imm    <="----------------";
					aRAout<="---";
					tellout<='0';
       end if; 
		 
		 if(WR_E='1') then 
               Iout <=Iin; 
               PCout<=PCin;
               opcode<=opcodein;
			     aluCout<=aluCin;
			     tellout<=tellin;
		         Imm    <=Immin;
					aRAout <=aRAin;
       end if;
  
		  
			 end if;
		end process;
end behave;